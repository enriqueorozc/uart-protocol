///////////////////////////////////////////////////////////////////////////////
// PROJECT: UART Communication System with Error Detection
///////////////////////////////////////////////////////////////////////////////
// AUTHORS: Enrique Orozco Jr. <enrique-orozco@outlook.com>
///////////////////////////////////////////////////////////////////////////////

module Uart_Receiver(uart_if uart);
endmodule