///////////////////////////////////////////////////////////////////////////////
// PROJECT: UART Communication System with Error Detection
///////////////////////////////////////////////////////////////////////////////
// AUTHORS: Enrique Orozco Jr. <enrique-orozco@outlook.com>
///////////////////////////////////////////////////////////////////////////////

module uart_rx(uart_if uart);
endmodule